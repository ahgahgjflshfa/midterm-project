`timescale 1ns/1ns
module TotalALU( clk, dataA, dataB, Signal, Output, reset );
    input reset ;
    input clk ;
    input [31:0] dataA ;
    input [31:0] dataB ;
    input [5:0] Signal ;
    output [31:0] Output ;

    //   Signal ( 6-bits)?
    //   AND  : 36
    //   OR   : 37
    //   ADD  : 32
    //   SUB  : 34
    //   SRL  : 2
    //   SLT  : 42
    //   MULTU : 25

    wire [31:0] temp ;

    parameter AND = 6'b100100;
    parameter OR  = 6'b100101;
    parameter ADD = 6'b100000;
    parameter SUB = 6'b100010;
    parameter SLT = 6'b101010;

    parameter SRL = 6'b000010;

    parameter MULTU = 6'd25;
    parameter MFHI = 6'b010000;
    parameter MFLO = 6'b010010;
    /*
    定義各種訊號
    */
    //============================
    wire carry;
    wire [5:0]  SignaltoALU ;
    wire [5:0]  SignaltoSHT ;
    wire [5:0]  SignaltoMUL ;
    wire [5:0]  SignaltoMUX ;
    wire [31:0] ALUOut, HiOut, LoOut, ShifterOut ;
    wire [31:0] dataOut ;
    wire [63:0] MULAns ;
    /*
    定義各種接線
    */
    //============================

    ALUControl ALUControl( .clk(clk), .Signal(Signal), .SignaltoALU(SignaltoALU), .SignaltoSHT(SignaltoSHT), .SignaltoMUL(SignaltoMUL), .SignaltoMUX(SignaltoMUX) );
    ALU ALU( .a(dataA), .b(dataB), .ctl(SignaltoALU), .result(ALUOut), .cin(0), .carry(carry));
    Multiplier Multiplier( .clk(clk), .dataA(dataA), .dataB(dataB), .Signal(SignaltoMUL), .dataOut(MULAns), .reset(reset) );
    Shifter Shifter( .a(dataA), .shamt(dataB), .Signal(SignaltoSHT), .result(ShifterOut));
    HiLo HiLo( .clk(clk), .MulAns(MulAns), .HiOut(HiOut), .LoOut(LoOut), .reset(reset));
    MUX MUX( .ALUOut(ALUOut), .HiOut(HiOut), .LoOut(LoOut), .Shifter(ShifterOut), .Signal(SignaltoMUX), .dataOut(dataOut) );
    /*
    建立各種module
    */
    assign Output = dataOut ;
endmodule