module Register_64bit();
    
endmodule