module tb();
    
endmodule