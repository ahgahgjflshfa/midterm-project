/*
    Title: 3 to 1 Mux
*/
module Mux_3to1(sel, in0, in1, in2);
endmodule